----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:23:54 12/02/2007 
-- Design Name: 
-- Module Name:    chargen - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity chargen is
	port (
		clk : in std_logic;
		output_addr : in std_logic_vector (11 downto 0);
		output_data : out std_logic_vector (3 downto 0)
	);
end chargen;

architecture Behavioral of chargen is
	signal oneSignal, zeroSignal : std_logic;
	signal xVector : std_logic_vector (3 downto 0);
begin
	oneSignal <= '1';
	zeroSignal <= '0';
	xVector <= "XXXX";
	
	RAMB16_S4_inst : RAMB16_S4 generic map (
		WRITE_MODE => "WRITE_FIRST",
		INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => X"9999999991111119911111199119911991199119911111199111111999999999",
		INIT_02 => X"aaaaaaaaa222222aa222222aa22aa22aa22aa22aa222222aa222222aaaaaaaaa",
		INIT_03 => X"bbbbbbbbb333333bb333333bb33bb33bb33bb33bb333333bb333333bbbbbbbbb",
		INIT_04 => X"ccccccccc444444cc444444cc44cc44cc44cc44cc444444cc444444ccccccccc",
		INIT_05 => X"ddddddddd555555dd555555dd55dd55dd55dd55dd555555dd555555ddddddddd",
		INIT_06 => X"eeeeeeeee666666ee666666ee66ee66ee66ee66ee666666ee666666eeeeeeeee",
		INIT_07 => X"fffffffff777777ff777777ff77ff77ff77ff77ff777777ff777777fffffffff",
		INIT_08 => X"7777777778888887788888877887788778877887788888877888888777777777",
		INIT_09 => X"2222222222222222222222222222222222222222222222222222222222222222",
		INIT_0a => X"2222222222222222222222227777777777777777222222222222222222222222",
		INIT_0b => X"2227722222277222222772222227722222277222222772222227722222277222",
		INIT_0c => X"2227722222277222227777227777777777777777227777222227722222277222",
		INIT_0d => X"2222222222222222222222227777222277777222227772222227722222277222",
		INIT_0e => X"2222222222222222222222222222777722277777222777222227722222277222",
		INIT_0f => X"2227722222277222227772227777722277772222222222222222222222222222",
		INIT_10 => X"2227722222277222222777222227777722227777222222222222222222222222",
		INIT_11 => X"0ef00ef00ef00ef00eeeeef00eeffef00ef00ef00eeeeef000ffff0000000000",
		INIT_12 => X"00eeeef00eeffef00ef00ef000effef00ef00ef00eeeeef000fffff000000000",
		INIT_13 => X"00eeee000efffef00ef00ef000000ef00ef00ef00eeeeef000ffff0000000000",
		INIT_14 => X"00eeeef00efffef00ef00ef00ef00ef00ef00ef00eeeeef000fffff000000000",
		INIT_15 => X"0eeeeef00ffffef000000ef000fffef000000ef00eeeeef00ffffff000000000",
		INIT_16 => X"00000ef000000ef000000ef000fffef000000ef00eeeeef00ffffff000000000",
		INIT_17 => X"00eeee000efffef00ef00ef00fff0ef000000ef00eeeeef000ffff0000000000",
		INIT_18 => X"0ef00ef00ef00ef00ef00ef00eeeeef00efffef00ef00ef00ef00ef000000000",
		INIT_19 => X"00eeef0000feef00000ef000000ef000000ef00000eeef0000ffff0000000000",
		INIT_1a => X"00eeee000eeffef00ef00ff00ef000000ef000000eeeeef00ffffff000000000",
		INIT_1b => X"0ee00ef00eee0ef000eeeef0000eeef000eefef00eef0ef00ff00ef000000000",
		INIT_1c => X"0eeeeef00ffffef000000ef000000ef000000ef000000ef000000ff000000000",
		INIT_1d => X"ee000ef0ee000ef0ee0e0ef0eeeeeef0eeefeef0eef0fef0ff000ff000000000",
		INIT_1e => X"ee000ef0eee00ef0eeee0ef0eefeeef0ef0feef0ef00fef0ff000ff000000000",
		INIT_1f => X"00eeee000eeffef00ef00ef00ef00ef00ef00ef00eeeeef000ffff0000000000",
		INIT_20 => X"00000ef000000ef000eeeef00eeffef00ee00ef00eeeeef000fffff000000000",
		INIT_21 => X"0eeeee000eeeeef00eef0ef00ee00ef00ee00ef00eeeeef000ffff0000000000",
		INIT_22 => X"0ee00ef000ee0ef000eeeef00eeffef00ee00ef00eeeeef000fffff000000000",
		INIT_23 => X"00eeeef00efffff00ef0000000ffff0000000ef00eeeeef00fffff0000000000",
		INIT_24 => X"000ef000000ef000000ef000000ef000000ef0000eeeeee00ffffff000000000",
		INIT_25 => X"00eeee000eeffef00ef00ef00ef00ef00ef00ef00ef00ef00ff00ff000000000",
		INIT_26 => X"000ef00000eeef0000eeef0000efff000ef00ef00ef00ef00ff00ff000000000",
		INIT_27 => X"0ee0ef00eefefef0ef0f0ef0ef0f0ef0ef000ef0ef000ef0ff000ff000000000",
		INIT_28 => X"ee000ef0eee0eef00eeeef0000eef0000eefef00eef0fef0ff000ff000000000",
		INIT_29 => X"000ef000000ef000000ef00000eeef000efffef00ef00ef00ff00ff000000000",
		INIT_2a => X"eeeeeef0fffeeef0000eef0000eef0000eef0000eeeeeef0fffffff000000000",
		INIT_2b => X"00eeee000eefeef00ef0eff00eeefef00eef0ef00eeeeef000ffff0000000000",
		INIT_2c => X"000ef000000ef000000ef000000ef000000eeef0000eef00000ff00000000000",
		INIT_2d => X"0eeeeef00ffeeef0000eef0000eef0000eef0ef00feeeef000ffff0000000000",
		INIT_2e => X"00eeee000eeffff00ff000f000eff0000ef000f00feeeef000ffff0000000000",
		INIT_2f => X"0ef000000ef000000ef000000eeeeef00eeffef00ef00ef00ff00ff000000000",
		INIT_30 => X"00eeeef00eeffff00ef0000000fffff0000000f00eeeeef00ffffff000000000",
		INIT_31 => X"00eeee000eeffef00ef00ef000fffef000000ef00feeeef000ffff0000000000",
		INIT_32 => X"0000ef000000ef00000eef0000eef0000eef00000eeeeef00ffffff000000000",
		INIT_33 => X"00eeee000eeffef00ef00ef000efff000ef00ef00eeeeef000ffff0000000000",
		INIT_34 => X"00eeee000eeffff00ef000000eeffe000ef00ef00eeeeef000ffff0000000000",
		INIT_35 => X"00000000000ef000000ff00000000000000ef000000ff0000000000000000000",
		INIT_36 => X"000ef000000ff00000000000000ef000000ef000000ef000000ff00000000000",
		INIT_37 => X"0000000000000000000000000eeeeef00ffffff0000000000000000000000000",
		INIT_38 => X"000ef000000ff000000000000000000000000000000000000000000000000000",
		INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3a => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3b => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3c => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3d => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3e => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3f => X"0000000000000000000000000000000000000000000000000000000000000000"
	) port map (
		DI => xVector,
		DO => output_data,
		ADDR => output_addr,
		CLK => clk,
		EN => oneSignal,
		SSR => zeroSignal,
		WE => zeroSignal
   );

end Behavioral;
